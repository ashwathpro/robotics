CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 82 1278 909
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 G:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 178 457 275
9961490 0
0
6 Title:
5 Name:
0
0
0
7
10 Capacitor~
219 544 436 0 1 5
0 0
0
0 0 832 90
3 1uF
11 0 32 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 0 0 0 0
1 C
5130 0 0
2
39777.3 0
0
10 Capacitor~
219 590 440 0 1 5
0 0
0
0 0 832 90
3 1uF
11 0 32 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 0 0 0 0
1 C
391 0 0
2
39777.3 0
0
7 Ground~
168 521 487 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3124 0 0
2
39777.3 0
0
9 Resistor~
219 620 337 0 1 5
0 0
0
0 0 864 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3421 0 0
2
39777.3 0
0
9 Resistor~
219 616 222 0 1 5
0 0
0
0 0 864 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8157 0 0
2
39777.3 0
0
2 +V
167 528 137 0 1 3
0 0
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5572 0 0
2
39777.3 0
0
10 555 Timer~
219 497 276 0 1 17
0 0
0
0 0 4928 0
3 555
-11 -36 10 -28
2 U1
-7 -46 7 -38
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
88 0 0 0 0 0 0 0
1 U
8901 0 0
2
39777.3 0
0
12
1 0 0 0 0 0 0 1 0 0 4 2
544 445
544 481
5 2 0 0 0 0 0 7 1 0 0 3
529 294
544 294
544 427
2 0 0 0 0 0 0 2 0 0 10 4
590 431
590 414
583 414
583 285
1 1 0 0 0 0 0 3 2 0 0 3
521 481
590 481
590 449
1 1 0 0 0 0 0 7 3 0 0 4
465 267
329 267
329 481
521 481
2 0 0 0 0 0 0 7 0 0 10 5
465 276
433 276
433 353
562 353
562 285
4 0 0 0 0 0 0 7 0 0 12 4
465 294
401 294
401 166
528 166
1 7 0 0 0 0 0 4 7 0 0 5
620 355
620 383
594 383
594 276
529 276
2 0 0 0 0 0 0 4 0 0 10 3
620 319
620 285
616 285
1 6 0 0 0 0 0 5 7 0 0 3
616 240
616 285
529 285
2 0 0 0 0 0 0 5 0 0 12 3
616 204
616 166
556 166
8 1 0 0 0 0 0 7 6 0 0 5
529 267
556 267
556 166
528 166
528 146
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
